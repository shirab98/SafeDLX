// Verilog test fixture created from schematic E:\adlx\B1\shirab2\Lab7\IO_SIMUL_VER\IO_SIM_DLX.sch - Thu Jan 09 16:09:19 2025

`timescale 1ns / 1ps

module IO_SIM_DLX_IO_SIM_DLX_sch_tb();

// Inputs
   reg STEP_IN;
   reg RESET_IN;
   reg CLK_IN;

// Output
   wire AS_N;
   wire [4:0] RD;
   wire IN_INIT;
   wire [11:0] STATE;
   wire STOP_N;
   wire WR_N;
	wire [31:0] PC;

// Bidirs

// Instantiate the UUT
   IO_SIM_DLX UUT (
		.AS_N(AS_N), 
		.RD(RD), 
		.IN_INIT(IN_INIT), 
		.STATE(STATE), 
		.STOP_N(STOP_N), 
		.STEP_IN(STEP_IN), 
		.WR_N(WR_N), 
		.RESET_IN(RESET_IN), 
		.CLK_IN(CLK_IN),
		.PC(PC)
   );
// Initialize Inputs
   
		initial 
		CLK_IN = 1;
		always 	 #10 CLK_IN = ~CLK_IN;
		initial begin
		#38;
      RESET_IN = 0;
		STEP_IN = 0 ;
		#80;
      RESET_IN = 1;
		#80;
		RESET_IN = 0;
		#80;
      STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		#80;
		STEP_IN = 0;
		#80;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
				STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		STEP_IN = 0;
		#160;
		STEP_IN = 1;
		#80;
		end
endmodule
