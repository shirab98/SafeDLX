library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity id is
Port ( id_num : out std_logic_vector(7 downto 0));
end id;

architecture Behavioral of id is

begin

   id_num <= X"4c";


end Behavioral;
