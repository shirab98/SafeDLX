`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:46:42 01/05/2025 
// Design Name: 
// Module Name:    DATA_COMPARATOR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DATA_COMPARATOR(
    input [31:0] S,
    input NEG,
    output COMP_OUT
    );

endmodule
